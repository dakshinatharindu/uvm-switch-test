package switch_pkg;

    // uvm
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // uvm_object
    `include "config_db.svh"

    // uvm_tests
    `include "switch_test.svh"
    
endpackage 